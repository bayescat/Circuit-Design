** Profile: "SCHEMATIC1-TRAN"  [ D:\OneDrive\OneDrive - Hyper Instrument\003_Simulation_Circuits\PSpice\TLV3501 Simulation\tlv3501-pspicefiles\schematic1\tran.sim ] 

** Creating circuit file "TRAN.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../TLV3501.lib" 
* From [PSPICE NETLIST] section of C:\Users\kimdo\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 500us 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
