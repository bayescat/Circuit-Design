** Profile: "SCHEMATIC1-tlv7011_sim"  [ D:\OneDrive\OneDrive - Hyper Instrument\003_Simulation_Circuits\OrCAD\TLV7011_Comparator Circuit\tlv7011-pspicefiles\schematic1\tlv7011_sim.sim ] 

** Creating circuit file "tlv7011_sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../tlv7011.lib" 
* From [PSPICE NETLIST] section of C:\Users\kimdo\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 2ms 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
