** Profile: "SCHEMATIC1-DITHER_RAS"  [ D:\OneDrive\OneDrive - Hyper Instrument\003_Simulation_Circuits\PSpice\RAS Circuit\dither_ras-pspicefiles\schematic1\dither_ras.sim ] 

** Creating circuit file "DITHER_RAS.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\kimdo\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 500ms 400ms 1 
.OPTIONS ADVCONV
.OPTIONS PIVTOL= 1.0E-12
.OPTIONS SOLVER= 0
.PROBE64 V(alias(*)) I(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
